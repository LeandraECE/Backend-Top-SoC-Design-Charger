##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Wed Dec 15 22:42:15 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERpower
  CLASS BLOCK ;
  SIZE 600.800000 BY 300.800000 ;
  FOREIGN BATCHARGERpower 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN iforcedbat
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 325.600000 300.160000 375.600000 300.800000 ;
      LAYER metal5 ;
        RECT 325.600000 300.160000 375.600000 300.800000 ;
    END
  END iforcedbat
  PIN vbatcurr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 200.520000 0.000000 200.680000 0.640000 ;
    END
  END vbatcurr
  PIN vsensbat
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 90.520000 0.000000 90.680000 0.640000 ;
    END
  END vsensbat
  PIN vref
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 100.520000 0.000000 100.680000 0.640000 ;
    END
  END vref
  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 0.000000 125.200000 0.640000 175.200000 ;
    END
  END vin
  PIN ibias1u
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 440.520000 0.000000 440.680000 0.640000 ;
    END
  END ibias1u
  PIN icc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 360.520000 0.000000 360.680000 0.640000 ;
    END
  END icc[7]
  PIN icc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 370.520000 0.000000 370.680000 0.640000 ;
    END
  END icc[6]
  PIN icc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 380.520000 0.000000 380.680000 0.640000 ;
    END
  END icc[5]
  PIN icc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 390.520000 0.000000 390.680000 0.640000 ;
    END
  END icc[4]
  PIN icc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 400.520000 0.000000 400.680000 0.640000 ;
    END
  END icc[3]
  PIN icc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 410.520000 0.000000 410.680000 0.640000 ;
    END
  END icc[2]
  PIN icc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 420.520000 0.000000 420.680000 0.640000 ;
    END
  END icc[1]
  PIN icc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 430.520000 0.000000 430.680000 0.640000 ;
    END
  END icc[0]
  PIN itc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 270.520000 0.000000 270.680000 0.640000 ;
    END
  END itc[7]
  PIN itc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 280.520000 0.000000 280.680000 0.640000 ;
    END
  END itc[6]
  PIN itc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 290.520000 0.000000 290.680000 0.640000 ;
    END
  END itc[5]
  PIN itc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 300.520000 0.000000 300.680000 0.640000 ;
    END
  END itc[4]
  PIN itc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 310.520000 0.000000 310.680000 0.640000 ;
    END
  END itc[3]
  PIN itc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 320.520000 0.000000 320.680000 0.640000 ;
    END
  END itc[2]
  PIN itc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 330.520000 0.000000 330.680000 0.640000 ;
    END
  END itc[1]
  PIN itc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 340.520000 0.000000 340.680000 0.640000 ;
    END
  END itc[0]
  PIN vcv[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 120.520000 0.000000 120.680000 0.640000 ;
    END
  END vcv[7]
  PIN vcv[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 130.520000 0.000000 130.680000 0.640000 ;
    END
  END vcv[6]
  PIN vcv[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 140.520000 0.000000 140.680000 0.640000 ;
    END
  END vcv[5]
  PIN vcv[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 150.520000 0.000000 150.680000 0.640000 ;
    END
  END vcv[4]
  PIN vcv[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 160.520000 0.000000 160.680000 0.640000 ;
    END
  END vcv[3]
  PIN vcv[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 170.520000 0.000000 170.680000 0.640000 ;
    END
  END vcv[2]
  PIN vcv[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 180.520000 0.000000 180.680000 0.640000 ;
    END
  END vcv[1]
  PIN vcv[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 190.520000 0.000000 190.680000 0.640000 ;
    END
  END vcv[0]
  PIN cc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 490.520000 0.000000 490.680000 0.640000 ;
    END
  END cc
  PIN tc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 210.520000 0.000000 210.680000 0.640000 ;
    END
  END tc
  PIN cv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 480.520000 0.000000 480.680000 0.640000 ;
    END
  END cv
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 450.520000 0.000000 450.680000 0.640000 ;
    END
  END en
  PIN sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 220.520000 0.000000 220.680000 0.640000 ;
    END
  END sel[3]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 230.520000 0.000000 230.680000 0.640000 ;
    END
  END sel[2]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 240.520000 0.000000 240.680000 0.640000 ;
    END
  END sel[1]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 250.520000 0.000000 250.680000 0.640000 ;
    END
  END sel[0]
  PIN avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 600.160000 160.100000 600.800000 161.100000 ;
    END
  END avdd
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 600.160000 119.300000 600.800000 120.300000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 600.160000 139.700000 600.800000 140.700000 ;
    END
  END dgnd
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 600.160000 180.500000 600.800000 181.500000 ;
    END
  END agnd
  PIN pgnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 0.100000 0.640000 1.100000 ;
    END
  END pgnd
  OBS
    LAYER metal1 ;
      RECT 0.000000 181.660000 600.800000 300.800000 ;
      RECT 0.000000 180.340000 600.000000 181.660000 ;
      RECT 0.000000 161.260000 600.800000 180.340000 ;
      RECT 0.000000 159.940000 600.000000 161.260000 ;
      RECT 0.000000 140.860000 600.800000 159.940000 ;
      RECT 0.000000 139.540000 600.000000 140.860000 ;
      RECT 0.000000 120.460000 600.800000 139.540000 ;
      RECT 0.000000 119.140000 600.000000 120.460000 ;
      RECT 0.000000 1.260000 600.800000 119.140000 ;
      RECT 0.800000 0.800000 600.800000 1.260000 ;
      RECT 490.840000 0.000000 600.800000 0.800000 ;
      RECT 480.840000 0.000000 490.360000 0.800000 ;
      RECT 450.840000 0.000000 480.360000 0.800000 ;
      RECT 440.840000 0.000000 450.360000 0.800000 ;
      RECT 430.840000 0.000000 440.360000 0.800000 ;
      RECT 420.840000 0.000000 430.360000 0.800000 ;
      RECT 410.840000 0.000000 420.360000 0.800000 ;
      RECT 400.840000 0.000000 410.360000 0.800000 ;
      RECT 390.840000 0.000000 400.360000 0.800000 ;
      RECT 380.840000 0.000000 390.360000 0.800000 ;
      RECT 370.840000 0.000000 380.360000 0.800000 ;
      RECT 360.840000 0.000000 370.360000 0.800000 ;
      RECT 340.840000 0.000000 360.360000 0.800000 ;
      RECT 330.840000 0.000000 340.360000 0.800000 ;
      RECT 320.840000 0.000000 330.360000 0.800000 ;
      RECT 310.840000 0.000000 320.360000 0.800000 ;
      RECT 300.840000 0.000000 310.360000 0.800000 ;
      RECT 290.840000 0.000000 300.360000 0.800000 ;
      RECT 280.840000 0.000000 290.360000 0.800000 ;
      RECT 270.840000 0.000000 280.360000 0.800000 ;
      RECT 250.840000 0.000000 270.360000 0.800000 ;
      RECT 240.840000 0.000000 250.360000 0.800000 ;
      RECT 230.840000 0.000000 240.360000 0.800000 ;
      RECT 220.840000 0.000000 230.360000 0.800000 ;
      RECT 210.840000 0.000000 220.360000 0.800000 ;
      RECT 200.840000 0.000000 210.360000 0.800000 ;
      RECT 190.840000 0.000000 200.360000 0.800000 ;
      RECT 180.840000 0.000000 190.360000 0.800000 ;
      RECT 170.840000 0.000000 180.360000 0.800000 ;
      RECT 160.840000 0.000000 170.360000 0.800000 ;
      RECT 150.840000 0.000000 160.360000 0.800000 ;
      RECT 140.840000 0.000000 150.360000 0.800000 ;
      RECT 130.840000 0.000000 140.360000 0.800000 ;
      RECT 120.840000 0.000000 130.360000 0.800000 ;
      RECT 100.840000 0.000000 120.360000 0.800000 ;
      RECT 90.840000 0.000000 100.360000 0.800000 ;
      RECT 0.800000 0.000000 90.360000 0.800000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 600.800000 300.800000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 600.800000 300.800000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 600.800000 300.800000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 600.800000 300.800000 ;
    LAYER metal6 ;
      RECT 375.880000 299.880000 600.800000 300.800000 ;
      RECT 0.000000 299.880000 325.320000 300.800000 ;
      RECT 0.000000 175.400000 600.800000 299.880000 ;
      RECT 0.840000 125.000000 600.800000 175.400000 ;
      RECT 0.000000 0.000000 600.800000 125.000000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 600.800000 300.800000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 600.800000 300.800000 ;
  END
END BATCHARGERpower

END LIBRARY
