##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Wed Jan  8 15:56:49 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERctr
  CLASS BLOCK ;
  SIZE 72.400000 BY 68.000000 ;
  FOREIGN BATCHARGERctr 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN cc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 71.880000 34.900000 72.400000 35.100000 ;
    END
  END cc
  PIN tc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 71.880000 34.100000 72.400000 34.300000 ;
    END
  END tc
  PIN cv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 71.880000 34.500000 72.400000 34.700000 ;
    END
  END cv
  PIN imonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 60.900000 0.000000 61.100000 0.520000 ;
    END
  END imonen
  PIN vmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 59.900000 0.000000 60.100000 0.520000 ;
    END
  END vmonen
  PIN tmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 61.900000 0.000000 62.100000 0.520000 ;
    END
  END tmonen
  PIN so
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 36.100000 67.480000 36.300000 68.000000 ;
    END
  END so
  PIN vbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 25.500000 0.000000 25.700000 0.520000 ;
    END
  END vbat[7]
  PIN vbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 24.700000 0.000000 24.900000 0.520000 ;
    END
  END vbat[6]
  PIN vbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 23.900000 0.000000 24.100000 0.520000 ;
    END
  END vbat[5]
  PIN vbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 23.100000 0.000000 23.300000 0.520000 ;
    END
  END vbat[4]
  PIN vbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 22.300000 0.000000 22.500000 0.520000 ;
    END
  END vbat[3]
  PIN vbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 21.500000 0.000000 21.700000 0.520000 ;
    END
  END vbat[2]
  PIN vbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 20.700000 0.000000 20.900000 0.520000 ;
    END
  END vbat[1]
  PIN vbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 19.900000 0.000000 20.100000 0.520000 ;
    END
  END vbat[0]
  PIN ibat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 38.900000 0.000000 39.100000 0.520000 ;
    END
  END ibat[7]
  PIN ibat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 38.100000 0.000000 38.300000 0.520000 ;
    END
  END ibat[6]
  PIN ibat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 37.300000 0.000000 37.500000 0.520000 ;
    END
  END ibat[5]
  PIN ibat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 36.500000 0.000000 36.700000 0.520000 ;
    END
  END ibat[4]
  PIN ibat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 35.700000 0.000000 35.900000 0.520000 ;
    END
  END ibat[3]
  PIN ibat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 34.900000 0.000000 35.100000 0.520000 ;
    END
  END ibat[2]
  PIN ibat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 34.100000 0.000000 34.300000 0.520000 ;
    END
  END ibat[1]
  PIN ibat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 33.300000 0.000000 33.500000 0.520000 ;
    END
  END ibat[0]
  PIN tbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 52.500000 0.000000 52.700000 0.520000 ;
    END
  END tbat[7]
  PIN tbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 51.700000 0.000000 51.900000 0.520000 ;
    END
  END tbat[6]
  PIN tbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 50.900000 0.000000 51.100000 0.520000 ;
    END
  END tbat[5]
  PIN tbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 50.100000 0.000000 50.300000 0.520000 ;
    END
  END tbat[4]
  PIN tbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 49.300000 0.000000 49.500000 0.520000 ;
    END
  END tbat[3]
  PIN tbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 48.500000 0.000000 48.700000 0.520000 ;
    END
  END tbat[2]
  PIN tbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 47.700000 0.000000 47.900000 0.520000 ;
    END
  END tbat[1]
  PIN tbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 46.900000 0.000000 47.100000 0.520000 ;
    END
  END tbat[0]
  PIN vcutoff[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 47.900000 0.520000 48.100000 ;
    END
  END vcutoff[7]
  PIN vcutoff[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 48.700000 0.520000 48.900000 ;
    END
  END vcutoff[6]
  PIN vcutoff[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 49.500000 0.520000 49.700000 ;
    END
  END vcutoff[5]
  PIN vcutoff[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 50.300000 0.520000 50.500000 ;
    END
  END vcutoff[4]
  PIN vcutoff[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 51.100000 0.520000 51.300000 ;
    END
  END vcutoff[3]
  PIN vcutoff[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 51.900000 0.520000 52.100000 ;
    END
  END vcutoff[2]
  PIN vcutoff[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 52.700000 0.520000 52.900000 ;
    END
  END vcutoff[1]
  PIN vcutoff[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 53.500000 0.520000 53.700000 ;
    END
  END vcutoff[0]
  PIN vpreset[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 41.500000 0.520000 41.700000 ;
    END
  END vpreset[7]
  PIN vpreset[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 42.300000 0.520000 42.500000 ;
    END
  END vpreset[6]
  PIN vpreset[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 43.100000 0.520000 43.300000 ;
    END
  END vpreset[5]
  PIN vpreset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 43.900000 0.520000 44.100000 ;
    END
  END vpreset[4]
  PIN vpreset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 44.700000 0.520000 44.900000 ;
    END
  END vpreset[3]
  PIN vpreset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 45.500000 0.520000 45.700000 ;
    END
  END vpreset[2]
  PIN vpreset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 46.300000 0.520000 46.500000 ;
    END
  END vpreset[1]
  PIN vpreset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 47.100000 0.520000 47.300000 ;
    END
  END vpreset[0]
  PIN tempmin[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 35.100000 0.520000 35.300000 ;
    END
  END tempmin[7]
  PIN tempmin[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 35.900000 0.520000 36.100000 ;
    END
  END tempmin[6]
  PIN tempmin[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 36.700000 0.520000 36.900000 ;
    END
  END tempmin[5]
  PIN tempmin[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 37.500000 0.520000 37.700000 ;
    END
  END tempmin[4]
  PIN tempmin[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 38.300000 0.520000 38.500000 ;
    END
  END tempmin[3]
  PIN tempmin[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 39.100000 0.520000 39.300000 ;
    END
  END tempmin[2]
  PIN tempmin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 39.900000 0.520000 40.100000 ;
    END
  END tempmin[1]
  PIN tempmin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 40.700000 0.520000 40.900000 ;
    END
  END tempmin[0]
  PIN tempmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 28.700000 0.520000 28.900000 ;
    END
  END tempmax[7]
  PIN tempmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 29.500000 0.520000 29.700000 ;
    END
  END tempmax[6]
  PIN tempmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 30.300000 0.520000 30.500000 ;
    END
  END tempmax[5]
  PIN tempmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 31.100000 0.520000 31.300000 ;
    END
  END tempmax[4]
  PIN tempmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 31.900000 0.520000 32.100000 ;
    END
  END tempmax[3]
  PIN tempmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 32.700000 0.520000 32.900000 ;
    END
  END tempmax[2]
  PIN tempmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 33.500000 0.520000 33.700000 ;
    END
  END tempmax[1]
  PIN tempmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 34.300000 0.520000 34.500000 ;
    END
  END tempmax[0]
  PIN tmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 22.300000 0.520000 22.500000 ;
    END
  END tmax[7]
  PIN tmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 23.100000 0.520000 23.300000 ;
    END
  END tmax[6]
  PIN tmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 23.900000 0.520000 24.100000 ;
    END
  END tmax[5]
  PIN tmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 24.700000 0.520000 24.900000 ;
    END
  END tmax[4]
  PIN tmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 25.500000 0.520000 25.700000 ;
    END
  END tmax[3]
  PIN tmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 26.300000 0.520000 26.500000 ;
    END
  END tmax[2]
  PIN tmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 27.100000 0.520000 27.300000 ;
    END
  END tmax[1]
  PIN tmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 27.900000 0.520000 28.100000 ;
    END
  END tmax[0]
  PIN iend[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 15.100000 0.520000 15.300000 ;
    END
  END iend[7]
  PIN iend[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 15.900000 0.520000 16.100000 ;
    END
  END iend[6]
  PIN iend[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 16.700000 0.520000 16.900000 ;
    END
  END iend[5]
  PIN iend[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 17.500000 0.520000 17.700000 ;
    END
  END iend[4]
  PIN iend[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 18.300000 0.520000 18.500000 ;
    END
  END iend[3]
  PIN iend[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 19.100000 0.520000 19.300000 ;
    END
  END iend[2]
  PIN iend[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 19.900000 0.520000 20.100000 ;
    END
  END iend[1]
  PIN iend[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 20.700000 0.520000 20.900000 ;
    END
  END iend[0]
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal4 ;
        RECT 9.900000 0.000000 10.100000 0.520000 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 10.700000 0.000000 10.900000 0.520000 ;
    END
  END en
  PIN rstz
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 11.500000 0.000000 11.700000 0.520000 ;
    END
  END rstz
  PIN vtok
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 21.500000 0.520000 21.700000 ;
    END
  END vtok
  PIN dvdd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
        RECT 11.900000 67.480000 12.100000 68.000000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
        RECT 9.900000 67.480000 10.100000 68.000000 ;
    END
  END dgnd
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 72.400000 68.000000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 72.400000 68.000000 ;
    LAYER metal3 ;
      RECT 0.000000 53.900000 72.400000 68.000000 ;
      RECT 0.720000 53.300000 72.400000 53.900000 ;
      RECT 0.000000 53.100000 72.400000 53.300000 ;
      RECT 0.720000 52.500000 72.400000 53.100000 ;
      RECT 0.000000 52.300000 72.400000 52.500000 ;
      RECT 0.720000 51.700000 72.400000 52.300000 ;
      RECT 0.000000 51.500000 72.400000 51.700000 ;
      RECT 0.720000 50.900000 72.400000 51.500000 ;
      RECT 0.000000 50.700000 72.400000 50.900000 ;
      RECT 0.720000 50.100000 72.400000 50.700000 ;
      RECT 0.000000 49.900000 72.400000 50.100000 ;
      RECT 0.720000 49.300000 72.400000 49.900000 ;
      RECT 0.000000 49.100000 72.400000 49.300000 ;
      RECT 0.720000 48.500000 72.400000 49.100000 ;
      RECT 0.000000 48.300000 72.400000 48.500000 ;
      RECT 0.720000 47.700000 72.400000 48.300000 ;
      RECT 0.000000 47.500000 72.400000 47.700000 ;
      RECT 0.720000 46.900000 72.400000 47.500000 ;
      RECT 0.000000 46.700000 72.400000 46.900000 ;
      RECT 0.720000 46.100000 72.400000 46.700000 ;
      RECT 0.000000 45.900000 72.400000 46.100000 ;
      RECT 0.720000 45.300000 72.400000 45.900000 ;
      RECT 0.000000 45.100000 72.400000 45.300000 ;
      RECT 0.720000 44.500000 72.400000 45.100000 ;
      RECT 0.000000 44.300000 72.400000 44.500000 ;
      RECT 0.720000 43.700000 72.400000 44.300000 ;
      RECT 0.000000 43.500000 72.400000 43.700000 ;
      RECT 0.720000 42.900000 72.400000 43.500000 ;
      RECT 0.000000 42.700000 72.400000 42.900000 ;
      RECT 0.720000 42.100000 72.400000 42.700000 ;
      RECT 0.000000 41.900000 72.400000 42.100000 ;
      RECT 0.720000 41.300000 72.400000 41.900000 ;
      RECT 0.000000 41.100000 72.400000 41.300000 ;
      RECT 0.720000 40.500000 72.400000 41.100000 ;
      RECT 0.000000 40.300000 72.400000 40.500000 ;
      RECT 0.720000 39.700000 72.400000 40.300000 ;
      RECT 0.000000 39.500000 72.400000 39.700000 ;
      RECT 0.720000 38.900000 72.400000 39.500000 ;
      RECT 0.000000 38.700000 72.400000 38.900000 ;
      RECT 0.720000 38.100000 72.400000 38.700000 ;
      RECT 0.000000 37.900000 72.400000 38.100000 ;
      RECT 0.720000 37.300000 72.400000 37.900000 ;
      RECT 0.000000 37.100000 72.400000 37.300000 ;
      RECT 0.720000 36.500000 72.400000 37.100000 ;
      RECT 0.000000 36.300000 72.400000 36.500000 ;
      RECT 0.720000 35.700000 72.400000 36.300000 ;
      RECT 0.000000 35.500000 72.400000 35.700000 ;
      RECT 0.720000 35.300000 72.400000 35.500000 ;
      RECT 0.720000 34.900000 71.680000 35.300000 ;
      RECT 0.000000 34.700000 71.680000 34.900000 ;
      RECT 0.720000 34.100000 71.680000 34.700000 ;
      RECT 0.000000 33.900000 71.680000 34.100000 ;
      RECT 0.720000 33.300000 72.400000 33.900000 ;
      RECT 0.000000 33.100000 72.400000 33.300000 ;
      RECT 0.720000 32.500000 72.400000 33.100000 ;
      RECT 0.000000 32.300000 72.400000 32.500000 ;
      RECT 0.720000 31.700000 72.400000 32.300000 ;
      RECT 0.000000 31.500000 72.400000 31.700000 ;
      RECT 0.720000 30.900000 72.400000 31.500000 ;
      RECT 0.000000 30.700000 72.400000 30.900000 ;
      RECT 0.720000 30.100000 72.400000 30.700000 ;
      RECT 0.000000 29.900000 72.400000 30.100000 ;
      RECT 0.720000 29.300000 72.400000 29.900000 ;
      RECT 0.000000 29.100000 72.400000 29.300000 ;
      RECT 0.720000 28.500000 72.400000 29.100000 ;
      RECT 0.000000 28.300000 72.400000 28.500000 ;
      RECT 0.720000 27.700000 72.400000 28.300000 ;
      RECT 0.000000 27.500000 72.400000 27.700000 ;
      RECT 0.720000 26.900000 72.400000 27.500000 ;
      RECT 0.000000 26.700000 72.400000 26.900000 ;
      RECT 0.720000 26.100000 72.400000 26.700000 ;
      RECT 0.000000 25.900000 72.400000 26.100000 ;
      RECT 0.720000 25.300000 72.400000 25.900000 ;
      RECT 0.000000 25.100000 72.400000 25.300000 ;
      RECT 0.720000 24.500000 72.400000 25.100000 ;
      RECT 0.000000 24.300000 72.400000 24.500000 ;
      RECT 0.720000 23.700000 72.400000 24.300000 ;
      RECT 0.000000 23.500000 72.400000 23.700000 ;
      RECT 0.720000 22.900000 72.400000 23.500000 ;
      RECT 0.000000 22.700000 72.400000 22.900000 ;
      RECT 0.720000 22.100000 72.400000 22.700000 ;
      RECT 0.000000 21.900000 72.400000 22.100000 ;
      RECT 0.720000 21.300000 72.400000 21.900000 ;
      RECT 0.000000 21.100000 72.400000 21.300000 ;
      RECT 0.720000 20.500000 72.400000 21.100000 ;
      RECT 0.000000 20.300000 72.400000 20.500000 ;
      RECT 0.720000 19.700000 72.400000 20.300000 ;
      RECT 0.000000 19.500000 72.400000 19.700000 ;
      RECT 0.720000 18.900000 72.400000 19.500000 ;
      RECT 0.000000 18.700000 72.400000 18.900000 ;
      RECT 0.720000 18.100000 72.400000 18.700000 ;
      RECT 0.000000 17.900000 72.400000 18.100000 ;
      RECT 0.720000 17.300000 72.400000 17.900000 ;
      RECT 0.000000 17.100000 72.400000 17.300000 ;
      RECT 0.720000 16.500000 72.400000 17.100000 ;
      RECT 0.000000 16.300000 72.400000 16.500000 ;
      RECT 0.720000 15.700000 72.400000 16.300000 ;
      RECT 0.000000 15.500000 72.400000 15.700000 ;
      RECT 0.720000 14.900000 72.400000 15.500000 ;
      RECT 0.000000 0.000000 72.400000 14.900000 ;
    LAYER metal4 ;
      RECT 36.500000 67.280000 72.400000 68.000000 ;
      RECT 12.300000 67.280000 35.900000 68.000000 ;
      RECT 10.300000 67.280000 11.700000 68.000000 ;
      RECT 0.000000 67.280000 9.700000 68.000000 ;
      RECT 0.000000 0.720000 72.400000 67.280000 ;
      RECT 62.300000 0.000000 72.400000 0.720000 ;
      RECT 61.300000 0.000000 61.700000 0.720000 ;
      RECT 60.300000 0.000000 60.700000 0.720000 ;
      RECT 52.900000 0.000000 59.700000 0.720000 ;
      RECT 52.100000 0.000000 52.300000 0.720000 ;
      RECT 51.300000 0.000000 51.500000 0.720000 ;
      RECT 50.500000 0.000000 50.700000 0.720000 ;
      RECT 49.700000 0.000000 49.900000 0.720000 ;
      RECT 48.900000 0.000000 49.100000 0.720000 ;
      RECT 48.100000 0.000000 48.300000 0.720000 ;
      RECT 47.300000 0.000000 47.500000 0.720000 ;
      RECT 39.300000 0.000000 46.700000 0.720000 ;
      RECT 38.500000 0.000000 38.700000 0.720000 ;
      RECT 37.700000 0.000000 37.900000 0.720000 ;
      RECT 36.900000 0.000000 37.100000 0.720000 ;
      RECT 36.100000 0.000000 36.300000 0.720000 ;
      RECT 35.300000 0.000000 35.500000 0.720000 ;
      RECT 34.500000 0.000000 34.700000 0.720000 ;
      RECT 33.700000 0.000000 33.900000 0.720000 ;
      RECT 25.900000 0.000000 33.100000 0.720000 ;
      RECT 25.100000 0.000000 25.300000 0.720000 ;
      RECT 24.300000 0.000000 24.500000 0.720000 ;
      RECT 23.500000 0.000000 23.700000 0.720000 ;
      RECT 22.700000 0.000000 22.900000 0.720000 ;
      RECT 21.900000 0.000000 22.100000 0.720000 ;
      RECT 21.100000 0.000000 21.300000 0.720000 ;
      RECT 20.300000 0.000000 20.500000 0.720000 ;
      RECT 11.900000 0.000000 19.700000 0.720000 ;
      RECT 11.100000 0.000000 11.300000 0.720000 ;
      RECT 10.300000 0.000000 10.500000 0.720000 ;
      RECT 0.000000 0.000000 9.700000 0.720000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 72.400000 68.000000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 72.400000 68.000000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 72.400000 68.000000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 72.400000 68.000000 ;
  END
END BATCHARGERctr

END LIBRARY
